library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ist_mem is
  port (
    clk, w : in std_logic;     
    pc     : in std_logic_vector(13 downto 0);
    addr_w : in std_logic_vector(13 downto 0);
    data   : in std_logic_vector(31 downto 0);
    ist    : out std_logic_vector(31 downto 0));
end ist_mem;

architecture behavior of ist_mem is

  -- moriya fib (register as displacement vesion)
  type ram_t is array (0 to 318) of std_logic_vector(31 downto 0);
  signal ram : ram_t := (x"00000000",
x"00000000",    
x"24400FF7",
x"24604268",
x"2C63000A",
x"2480000A",
x"74400003",
x"6C820000",
x"D00000CF",
x"04A02000",
x"64820000",
x"6CA20001",
x"6C820000",
x"D00000BC",
x"64A20000",
x"64C20001",
x"6C820002",
x"6CC20001",
x"6CA20000",
x"04802800",
x"04A03000",
x"D00000BC",
x"64A20000",
x"64C20001",
x"6C820003",
x"04802800",
x"04A03000",
x"D00000BC",
x"64A20002",
x"6C820004",
x"04802800",
x"D00000EF",
x"64A20003",
x"6C820005",
x"04802800",
x"D00000EF",
x"64A20004",
x"6C820006",
x"04802800",
x"D00000EF",
x"04C02000",
x"24800000",
x"64A20005",
x"04852000",
x"64840000",
x"24E00000",
x"74400002",
x"04843800",
x"7C440000",
x"24800000",
x"04852000",
x"64840000",
x"24E00001",
x"74400003",
x"04843800",
x"7C440000",
x"24800000",
x"04852000",
x"64840000",
x"24E00002",
x"74400003",
x"04843800",
x"7C440000",
x"24800001",
x"04852000",
x"64840000",
x"24E00000",
x"74400003",
x"04843800",
x"7C440000",
x"24800001",
x"04852000",
x"64840000",
x"24E00001",
x"74400001",
x"04843800",
x"7C440000",
x"24800001",
x"04852000",
x"64840000",
x"24E00002",
x"74400003",
x"04843800",
x"7C440000",
x"24800002",
x"04852000",
x"64840000",
x"24E00000",
x"74400003",
x"04843800",
x"7C440000",
x"24800002",
x"04852000",
x"64840000",
x"24E00001",
x"74400003",
x"04843800",
x"7C440000",
x"24800002",
x"04852000",
x"64840000",
x"24E00002",
x"74400000",
x"04843800",
x"7C440000",
x"24800000",
x"64E20006",
x"04872000",
x"64840000",
x"25000000",
x"74400002",
x"04844000",
x"7C440000",
x"24800000",
x"04872000",
x"64840000",
x"25000001",
x"74400003",
x"04844000",
x"7C440000",
x"24800000",
x"04872000",
x"64840000",
x"25000002",
x"74400003",
x"04844000",
x"7C440000",
x"24800001",
x"04872000",
x"64840000",
x"25000000",
x"74400003",
x"04844000",
x"7C440000",
x"24800001",
x"04872000",
x"64840000",
x"25000001",
x"74400001",
x"04844000",
x"7C440000",
x"24800001",
x"04872000",
x"64840000",
x"25000002",
x"74400003",
x"04844000",
x"7C440000",
x"24800002",
x"04872000",
x"64840000",
x"25000000",
x"74400003",
x"04844000",
x"7C440000",
x"24800002",
x"04872000",
x"64840000",
x"25000001",
x"74400003",
x"04844000",
x"7C440000",
x"24800002",
x"04872000",
x"64840000",
x"25000002",
x"74400000",
x"04844000",
x"7C440000",
x"6CC20007",
x"04802800",
x"04A03800",
x"D0000134",
x"24800002",
x"64A20007",
x"04852000",
x"64840000",
x"24A00002",
x"04842800",
x"74440000",
x"D0000136",
x"C0000139",
x"84A00002",
x"E0000000",
x"7C440000",
x"28A50001",
x"24840001",
x"C00000B6",
x"28420001",
x"04C01800",
x"04632000",
x"6CC20000",
x"04203000",
x"04C02800",
x"04A02000",
x"04800800",
x"D00000C9",
x"64820000",
x"04802000",
x"24420001",
x"E0000000",
x"84A00002",
x"E0000000",
x"6CC40000",
x"28A50001",
x"24840001",
x"C00000C9",
x"28420001",
x"04A01800",
x"04632000",
x"6CA20000",
x"04202800",
x"04A02000",
x"04800800",
x"D00000B6",
x"64820000",
x"04802000",
x"24420001",
x"E0000000",
x"28420002",
x"24C0000A",
x"84A60004",
x"04802000",
x"24420002",
x"E0000000",
x"74400003",
x"6CA20000",
x"6C820001",
x"04803000",
x"D00000CF",
x"64A20000",
x"64C20001",
x"04E62800",
x"6C870000",
x"24800001",
x"04A52000",
x"04803000",
x"24420002",
x"C00000DB",
x"24A00000",
x"C00000DB",
x"2540000A",
x"850A0002",
x"E0000000",
x"05463800",
x"654A0000",
x"05663800",
x"656B0000",
x"056B4800",
x"744B0000",
x"05643800",
x"656B0000",
x"056B4000",
x"746B0000",
x"05654000",
x"656B0000",
x"056B4800",
x"748B0000",
x"48632000",
x"40421800",
x"054A4800",
x"7C4A0000",
x"25400001",
x"05085000",
x"C00000F1",
x"28420005",
x"2520000A",
x"85090003",
x"24420005",
x"E0000000",
x"25200000",
x"6CE20000",
x"6CC20001",
x"6CA20002",
x"6C820003",
x"6D020004",
x"04204800",
x"05204000",
x"05000800",
x"D00000F1",
x"24800001",
x"64A20004",
x"05052000",
x"64820003",
x"64A20002",
x"64C20001",
x"64E20000",
x"24420005",
x"C0000109",
x"28420004",
x"2500000A",
x"84E80003",
x"24420004",
x"E0000000",
x"25000000",
x"6CC20000",
x"6CA20001",
x"6C820002",
x"6CE20003",
x"D0000109",
x"24800001",
x"64A20003",
x"04E52000",
x"64820002",
x"64A20001",
x"64C20000",
x"24420004",
x"C0000121",
x"24E00000",
x"C0000121",
x"74600003",
x"40421800",
x"E0000000",
x"6C800FFF",
x"40420000",
x"C000013A",
x"00000000",
x"00000000",
x"FFFFFFFF");
                           
begin

  write: process(clk)
  begin
    if rising_edge(clk) then
      ist <= ram(conv_integer(pc(8 downto 0)));
      if w = '1' then
        ram(conv_integer(addr_w)) <= data;
      end if;
    end if;
  end process;
  
end behavior;
    
